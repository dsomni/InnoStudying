module ex2(i1,i2,b0,a,b,c,d,e,f,d4,d6,d8,d10,d12,d14);
	input i1,i2;
	output b0,a,b,c,d,e,f,d4,d6,d8,d10,d12,d14;
	
	assign b0 = i1;
	assign a = i1;
	assign b = i1;
	assign c = i1;
	assign d = i1;
	assign e = i1;
	assign f = i1;
	
	assign d4 = i2;
	assign d6 = i2;
	assign d8 = i2;
	assign d10 = i2;
	assign d12 = i2;
	assign d14 = i2;
	
endmodule
	
	