module ex3(i1, b0, b1,b2, b3, b4, b5, b6,b7,a);
	input i1;
	output b0, b1,b2, b3, b4, b5, b6,b7,a;
	
	assign b0 = i1;
	assign b1 = i1;
   assign b2 = i1;
	assign b3 = i1;
	assign b4 = i1;
	assign b5 = i1;
	assign b6 = i1;
	assign b7 = i1;
	assign a = 0;


endmodule